library IEEE;
use IEEE.STD_LOGIC_1164.all;

package defines is
  constant directory : string := "F:\HDL\Synthesizer\repo\Oscillator_2.0\src\";
  
end package defines;